module not_gate_df(a,y);
input a;
output wire y;
assign y = ~a;
endmodule
