module nor_gate(a,b,y);
input a,b;
output wire y;
nor(y,a,b);
endmodule
