module xor_gate(a,b,y);
input a,b;
output wire y;
xor(y,a,b);
endmodule
