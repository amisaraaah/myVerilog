module not_gate(a,y);
input a;
output wire y;
not(y,a);
endmodule
