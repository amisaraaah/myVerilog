module xnor_gate(a,b,y);
input a,b;
output wire y;
xnor(y,a,b);
endmodule
