module and_gate(a,b,y);
input a,b;
output wire y;
and(y,a,b);
endmodule
