module or_gate(a,b,y);
input a,b;
output wire y;
or(y,a,b);
endmodule